@00000000
01 10 04 00 10 00 2E 22 02 32 02 42 02 52 02 62 
82 01 83 01 84 01 85 01 86 01 09 60 04 00 00 00 
08 70 04 00 00 00 1A 00 00 00 10 10 0F 00 0F 00 
