@00000000
2E 22 2E 33 2E 44 2E 55 2E 66 82 01 83 01 84 01 
85 01 86 01 82 01 83 01 84 01 85 01 86 01 82 01 
83 01 84 01 85 01 86 01 
