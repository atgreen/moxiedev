// cpu_ififo.v - The instruction FIFO unit
//
// Copyright (c) 2010, 2011 Anthony Green.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
// 
// The above named program is free software; you can redistribute it
// and/or modify it under the terms of the GNU General Public License
// version 2 as published by the Free Software Foundation.
// 
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty
// of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA
// 02110-1301, USA.

module cpu_ififo (/*AUTOARG*/
  // Outputs
  opcode_o, operand_o, valid_o, empty_o, full_o,
  // Inputs
  rst_i, clk_i, write_en_i, read_en_i, data_i
  );
  
  // --- Clock and Reset ------------------------------------------
  input  rst_i, clk_i;

  input write_en_i ; // assert high to write data
  input read_en_i ; // assert high to read data

  input [31:0] data_i ; // data to write
  
  output [15:0] opcode_o; // opcode_o for newly read instruction
  output [31:0] operand_o; // data operand_o for newly read instruction
  output [0:0]	valid_o;
  output [0:0]	empty_o ;
  output [0:0]	full_o ;
  
  reg [1:0]    read_ptr, write_ptr; // write and read pointers
  reg [2:0]    ptr_gap; // gap between the pointers
  reg [15:0]   opcode_o;
  reg [31:0]   operand_o;
  reg [0:0]    valid_o;
  reg [0:0]    full_o;
  reg [15:0]   buffer[3:0]; // instruction buffer

  wire [0:0]   can_write_32, can_read_16, can_read_48;
  wire [0:0]   buffer_full,  buffer_empty;
  
  assign can_write_32 = ((ptr_gap == 0) || (ptr_gap == 1) || (ptr_gap == 2));
  assign can_read_16 = (ptr_gap != 0);
  assign can_read_48 =  ((ptr_gap != 0) && (ptr_gap != 1) && (ptr_gap != 2));
  assign buffer_full = ptr_gap == 4;
  assign buffer_empty = ptr_gap == 0;

  assign empty_o = buffer_empty;

  // This is a rediculous bit of logic.  We should try to recode the
  // moxie instructions so that we can determine the length with less
  // logic.
  function [0:0] is_long_insn;
    input [7:0] op;
    is_long_insn = ((op == 8'h01) //  ldi.l
		    || (op == 8'h03) // jsra
		    || (op == 8'h08) // lda.l
		    || (op == 8'h09) // sta.l
		    || (op == 8'h0c) // ldo.l
		    || (op == 8'h0d) // sto.l
		    || (op == 8'h1a) // jmpa
		    || (op == 8'h1b) // ldi.b
		    || (op == 8'h1d) // lda.b
		    || (op == 8'h1f) // sta.b
		    || (op == 8'h20) // ldi.s
		    || (op == 8'h22) // lda.s
		    || (op == 8'h24) // sta.s
		    || (op == 8'h25) // jmp
		    || (op == 8'h30) // swi
		    || (op == 8'h36) // ldo.b
		    || (op == 8'h37) // sto.b
		    || (op == 8'h38) // ldo.s
		    || (op == 8'h39) // sto.s
		    // Easy optimization.. all insns with two high bits on
		    // are 48-bits long.
		    || (op == 8'hc0) // beq
		    || (op == 8'hc4) // bne
		    || (op == 8'hc8) // blt
		    || (op == 8'hcc) // bgt
		    || (op == 8'hd0) // bltu
		    || (op == 8'hd4) // bgtu
		    || (op == 8'hd8) // bge
		    || (op == 8'hdc) // ble
		    || (op == 8'he0) // bgeu
		    || (op == 8'he4)); // bleu
  endfunction

  always @(posedge clk_i or posedge rst_i)
    if (rst_i == 1) begin
      opcode_o <= 0;
      operand_o <= 0;
      read_ptr <= 0;
      write_ptr <= 0;
      ptr_gap <= 0;
      full_o <= 0;
      valid_o <= 0;
    end else begin
      // $display ("A %x buffer[read_ptr] = 0x%x", read_ptr, buffer[read_ptr][15:8]);
      // $display ("A BUFFER = 0x%x%x%x%x", buffer[0], buffer[1], buffer[2], buffer[3]);
      // $display ("A buffer_empty = %x", buffer_empty);
      // $display ("A ptr_gap = 0x%x", ptr_gap);
      // $display ("A 0x%x", !is_long_insn(buffer[read_ptr][15:8]));
      // $display ("A 0x%x", buffer[read_ptr][15:8]);
      if (buffer_empty ? !is_long_insn(data_i[31:24]) : !is_long_insn(buffer[read_ptr][15:8])) begin
	// This is a 16-bit instruction (either from input or from buffer).
	//	$display ("B");
	if (write_en_i && (!read_en_i) && (can_write_32)) begin
	  //	  $display ("Z");
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[(write_ptr+1)%4] <= data_i[15:0];
	  write_ptr <= (write_ptr + 2) % 4;
	  valid_o <= 0;
	  ptr_gap = ptr_gap + 2;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if ((!write_en_i) && read_en_i && (can_read_16)) begin
	  // $display ("Y");
	  opcode_o <= buffer[read_ptr];
	  valid_o <= 1;
	  read_ptr <= (read_ptr + 1) % 4;
	  ptr_gap = ptr_gap - 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if (write_en_i && read_en_i && buffer_empty) begin
	  //	   $display ("X");
	  opcode_o <= data_i[31:16];
	  buffer[0] <= data_i[15:0];
	  write_ptr <= 1;
	  read_ptr <= 0;
	  ptr_gap = 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  valid_o <= 1;
	end
	else if (write_en_i && read_en_i && buffer_full) begin
	  //	   $display ("W- ERROR");
	  opcode_o <= buffer[read_ptr];
	  valid_o <= 1;
	  read_ptr <= (read_ptr + 1) % 4;
	  ptr_gap = ptr_gap - 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if (write_en_i && read_en_i && (can_write_32) && (can_read_16)) begin
	  //	   $display ("V");
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[(write_ptr+1)%4] <= data_i[15:0];
	  write_ptr <= (write_ptr + 2) % 4;
	  opcode_o <= buffer[read_ptr];
	  read_ptr <= (read_ptr + 1) % 4;
	  valid_o <= 1;
	  ptr_gap = ptr_gap + 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  // #1 $display ("V - %x %x %x %x %x %x", write_en_i, read_en_i, write_ptr, read_ptr, ptr_gap, 
//		       full_o);
	end 
	else begin
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  // #1 $display ("U - ERROR %x %x %x %x %x %x", write_en_i, read_en_i, write_ptr, read_ptr, ptr
	  // _gap, full_o);
	end
      end else begin
	// $display ("C w %x r %x w32 %x", write_en_i, read_en_i, can_write_32);
	if (write_en_i && (!read_en_i) && (can_write_32)) begin
	  //	   $display ("D");
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[write_ptr+1] <= data_i[15:0];
	  write_ptr <= write_ptr + 2;
	  ptr_gap = ptr_gap + 2;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if ((!write_en_i) && read_en_i && (can_read_48)) begin
	  //	   $display ("E");
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= buffer[read_ptr+1];
	  operand_o[15:0] <= buffer[read_ptr+2];
	  valid_o <= 1;
	  read_ptr <= read_ptr + 3;
	  ptr_gap = ptr_gap - 3;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  //	  #1 $display ("eee... opcode_o = %x, %x", opcode_o, is_long_insn(opcode_o));
	  //	  #1 $display ("eee... buffer = 0x%x%x%x%x", buffer[read_ptr], buffer[read_ptr+1], buffer[read_ptr+2], buffer[read_ptr+3]);
	end
	else if (write_en_i && read_en_i && buffer_empty) begin
	  //	   $display ("F data = 0x%x", data_i);
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[write_ptr+1] <= data_i[15:0];
	  write_ptr <= write_ptr + 2;
	  valid_o <= 0;
	  ptr_gap = ptr_gap + 2;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  //	  // #1 $display ("f... buffer = 0x%x%x%x%x", buffer[read_ptr], buffer[read_ptr+1], buffer[read_
	    // ptr+2], buffer[read_ptr+3]);
	end
	else if (write_en_i && read_en_i && buffer_full) begin
	  //	   $display ("G");
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= buffer[read_ptr+1];
	  operand_o[15:0] <= buffer[read_ptr+2];
	  valid_o <= 1;
	  read_ptr <= read_ptr + 3;
	  ptr_gap = ptr_gap - 3;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if (write_en_i && read_en_i && (can_write_32) && (can_read_48)) begin
	  //	   $display ("H");
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[write_ptr+1] <= data_i[15:0];
	  write_ptr <= write_ptr + 2;
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= buffer[read_ptr+1];
	  operand_o[15:0] <= buffer[read_ptr+2];
	  read_ptr <= read_ptr + 3;
	  valid_o <= 1;
	  ptr_gap = ptr_gap - 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	end
	else if (write_en_i && read_en_i && (ptr_gap == 2)) begin
	  //	   $display ("I");
	  buffer[(write_ptr)%4] <= data_i[31:16];
	  buffer[(write_ptr+1)%4] <= data_i[15:0];
	  write_ptr <= (write_ptr + 2) % 4;
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= buffer[(read_ptr+1)%4];
	  operand_o[15:0] <= data_i[31:16];
	  read_ptr <= (read_ptr + 3) % 4;
	  valid_o <= 1;
	  ptr_gap = 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  // #1 $display ("opcode = 0x%x, operand = 0x%x, valid = %x", opcode_o, operand_o, valid_o );
	  // #1 $display ("i... rbuffer[0x%x] = 0x%x%x%x%x", read_ptr, buffer[read_ptr], buffer[(read_ptr+1)%4], buffer[(read_ptr+2)%4], buffer[(read_ptr+3)%4]);
	  // #1 $display ("i... wbuffer[0x%x] = 0x%x%x%x%x", write_ptr, buffer[write_ptr], buffer[(write_ptr+1)%4], buffer[(write_ptr+2)%4], buffer[(write_ptr+3)%4]);
	  // #1 $display ("0x%x 0x%x 0x%x 0x%x", write_ptr, write_ptr+1, write_ptr+2, write_ptr+3);
	end
	else if (write_en_i && read_en_i && (ptr_gap == 1)) begin
	  //	  $display ("J data = 0x%x, read_ptr = 0x%x", data_i, read_ptr);
	  //	  $display ("i... rbuffer[0x%x] = 0x%x%x%x%x", read_ptr, buffer[read_ptr], buffer[(read_ptr+1)%4], buffer[(read_ptr+2)%4], buffer[(read_ptr+3)%4]);
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= data_i[31:16];
	  operand_o[15:0] <= data_i[15:0];
	  read_ptr <= (read_ptr + 1) % 4;
	  valid_o <= 1;
	  ptr_gap = 0;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  // #1 $display ("j... buffer[0x%x] = 0x%x%x%x%x", read_ptr, buffer[read_ptr], buffer[(read_ptr
	  //	    +1)%4], buffer[(read_ptr+2)%4], buffer[(read_ptr+3)%4]);
	end 
	else if (write_en_i && read_en_i && (ptr_gap == 3)) begin
	  //	   $display ("K data = 0x%x", data_i);
	  buffer[write_ptr] <= data_i[31:16];
	  buffer[write_ptr+1] <= data_i[15:0];
	  write_ptr <= write_ptr + 2;
	  opcode_o <= buffer[read_ptr];
	  operand_o[31:16] <= buffer[(read_ptr+1)%4];
	  operand_o[15:0] <= buffer[(read_ptr+2)%4];
	  read_ptr <= read_ptr + 3;
	  valid_o <= 1;
	  ptr_gap = ptr_gap - 1;
	  full_o = ((ptr_gap == 3) || (ptr_gap == 4));
	  // #1 $display ("k... buffer[0x%x] = 0x%x%x%x%x", read_ptr, buffer[read_ptr], buffer[(read_ptr
	  // +1)%4], buffer[(read_ptr+2)%4], buffer[(read_ptr+3)%4]);
	end 
	  // else #1 $display ("L ERROR ptr_gap = 0x%x", ptr_gap);
      end  
    end
endmodule

