@00001000
01 10 00 40 00 00 01 00 00 00 00 00 91 0C 01 20 
00 00 53 84 01 30 00 00 53 C4 29 32 0D 13 00 00 
00 08 01 30 00 00 00 00 03 00 00 00 11 6C 81 0C 
03 00 00 00 49 FE 01 20 00 00 4A 0C 03 00 00 00 
11 22 08 20 00 00 00 04 01 30 00 00 00 08 03 00 
00 00 11 0C 03 00 00 00 11 38 06 18 06 19 06 1A 
06 1B 91 18 01 30 00 00 00 18 1D 20 00 00 53 84 
28 23 27 23 01 30 00 00 00 00 0E 23 C4 26 08 20 
00 00 53 88 01 80 00 00 53 7C 01 90 00 00 53 78 
29 89 01 A0 00 00 00 02 2D 8A 98 01 0E 28 E0 0F 
82 01 09 20 00 00 53 88 28 2A 02 39 05 32 0A 23 
19 20 08 20 00 00 53 88 0E 28 D3 F3 1B 20 00 00 
00 01 1F 20 00 00 53 84 02 70 97 10 07 7B 07 7A 
07 79 07 78 04 00 91 18 04 00 06 1B 91 18 01 20 
00 00 00 00 08 30 00 00 53 80 0E 32 C0 0A 01 30 
00 00 00 00 0E 32 C0 05 01 20 00 00 53 80 19 30 
02 70 97 04 07 7B 04 00 91 18 04 00 91 18 01 20 
00 00 4A 14 03 00 00 00 13 6C 01 20 00 00 00 00 
04 00 91 18 02 32 01 20 00 00 00 00 02 42 02 52 
03 00 00 00 14 2E 04 00 06 18 06 1B 91 18 02 82 
01 30 00 00 00 00 03 00 00 00 15 82 08 20 00 00 
4A 24 0C 32 00 00 00 3C 01 40 00 00 00 00 0E 34 
C0 02 19 30 02 28 03 00 00 00 49 E0 06 18 06 19 
06 1A 06 1B 02 52 01 E0 00 00 00 03 02 82 26 8E 
01 60 00 00 00 00 0E 86 C0 11 0E 46 C0 78 94 01 
02 83 1A 00 00 00 11 9E 0E 46 C0 71 94 01 1E 58 
85 01 02 95 26 9E 0E 96 C7 F8 01 60 00 00 00 03 
0E 46 E4 5A 01 90 00 00 00 FF 02 63 26 69 02 96 
02 65 01 80 00 00 00 08 02 A9 28 A8 02 8A 2B 89 
01 E0 00 00 00 10 02 98 28 9E 02 E9 2B E8 01 90 
00 00 00 0F 0E 49 E4 24 02 65 02 84 0B 6E 0D 6E 
00 00 00 04 0D 6E 00 00 00 08 0D 6E 00 00 00 0C 
86 10 98 10 0E 89 D7 F3 94 10 01 80 00 00 00 04 
02 64 27 68 86 01 28 68 05 56 02 65 01 50 00 00 
00 0F 26 45 01 50 00 00 00 03 0E 45 E4 1C 01 50 
00 00 00 00 01 80 00 00 00 03 02 96 05 95 0B 9E 
85 04 02 94 29 95 0E 98 D7 F9 94 04 01 80 00 00 
00 02 02 54 27 58 85 01 28 58 05 65 01 50 00 00 
00 03 26 45 02 56 01 60 00 00 00 00 0E 46 C0 07 
02 85 05 86 1E 83 86 01 0E 46 C7 FB 02 70 97 10 
07 7B 07 7A 07 79 07 78 04 00 06 18 06 19 06 1B 
91 34 02 82 02 93 02 23 03 00 00 00 13 7E 0D 09 
FF FF FF D8 0D 02 FF FF FF DC 01 30 00 00 4A 2C 
0D 03 FF FF FF E0 01 30 00 00 00 01 0D 03 FF FF 
FF E4 05 23 0D 02 FF FF FF F0 02 20 92 28 0D 02 
FF FF FF E8 01 20 00 00 00 02 0D 02 FF FF FF EC 
08 20 00 00 4B 34 0C 22 00 00 00 08 38 42 00 00 
00 0C 01 30 00 00 00 10 02 54 28 53 27 53 01 30 
00 00 20 00 26 53 01 60 00 00 00 00 0E 56 C4 0F 
2B 43 39 24 00 00 00 0C 0C 32 00 00 00 64 01 40 
FF FF DF FF 26 34 0D 23 00 00 00 64 02 28 0C 38 
00 00 00 08 02 40 94 18 03 00 00 00 17 5E 01 30 
00 00 00 00 0E 23 C4 0A 01 20 00 00 00 0A 02 70 
97 0C 07 7B 07 79 07 78 04 00 01 20 FF FF FF FF 
02 70 97 0C 07 7B 07 79 07 78 04 00 91 18 02 32 
08 20 00 00 4B 34 03 00 00 00 12 8A 04 00 06 18 
06 1B 01 60 00 00 00 03 02 32 26 36 01 40 00 00 
00 00 0E 34 C0 49 01 50 00 00 00 18 1C 32 28 35 
2D 35 0E 34 C0 3B 02 32 1A 00 00 00 13 B8 1C E3 
28 E5 2D E5 0E E4 C0 31 83 01 02 E3 26 E6 0E E4 
C7 F7 0A 53 01 60 FE FE FE FF 02 45 05 46 2C 55 
26 45 01 50 80 80 80 80 26 45 01 80 00 00 00 00 
0E 48 C4 0A 83 04 0A 83 02 E8 05 E6 2C 88 26 E8 
26 E5 0E E4 C3 F8 01 40 00 00 00 18 1C 63 28 64 
2D 64 01 50 00 00 00 00 0E 65 C0 07 83 01 1C 63 
28 64 2D 64 0E 65 C7 FB 29 32 02 23 02 70 97 08 
07 7B 07 78 04 00 02 32 1A 00 00 00 13 C2 06 18 
06 19 06 1A 06 1B 91 24 02 82 08 90 00 00 4A 24 
0C 29 00 00 01 48 01 60 00 00 00 00 0E 26 C0 52 
0C A2 00 00 00 04 01 60 00 00 00 1F 0E A6 CC 56 
02 6A 86 01 01 90 00 00 00 00 0E 89 C4 16 8A 02 
01 40 00 00 00 02 28 A4 02 42 05 4A 0B 43 0D 26 
00 00 00 04 01 20 00 00 00 00 02 70 97 10 07 7B 
07 7A 07 79 07 78 04 00 02 9A 89 22 01 60 00 00 
00 02 28 96 02 B2 05 B9 0B B4 01 40 00 00 00 01 
28 4A 0C 92 00 00 01 88 2B 94 0D 29 00 00 01 88 
02 9A 89 42 28 96 02 B2 05 B9 0B B5 0E 86 C0 06 
02 6A 86 01 1A 00 00 00 14 6E 0C 52 00 00 01 8C 
2B 54 0D 25 00 00 01 8C 02 6A 86 01 1A 00 00 00 
14 6E 01 20 00 00 01 4C 02 69 05 62 02 26 0D 96 
00 00 01 48 1A 00 00 00 14 50 01 60 00 00 00 00 
01 A0 00 00 00 00 0E 6A C4 07 01 20 FF FF FF FF 
1A 00 00 00 14 8A 01 20 00 00 01 90 0D 03 FF FF 
FF EC 0D 04 FF FF FF E8 0D 05 FF FF FF E4 19 60 
0E 2A 0C 30 FF FF FF EC 0C 40 FF FF FF E8 0C 50 
FF FF FF E4 C3 E3 0D 2A 00 00 00 04 0C 69 00 00 
01 48 0B 26 0D 92 00 00 01 48 0D 2A 00 00 01 88 
0D 2A 00 00 01 8C 01 60 00 00 00 01 1A 00 00 00 
14 64 06 18 06 19 06 1A 06 1B 06 1C 06 1D 91 28 
0D 02 00 00 00 0C 02 43 01 90 00 00 00 00 01 20 
00 00 01 48 08 30 00 00 4A 24 05 32 0D 03 FF FF 
FF E4 08 20 00 00 4A 24 0C D2 00 00 01 48 0E D9 
C0 2A 0C 60 FF FF FF E4 0C CD 00 00 00 04 02 8C 
98 01 0E 89 C8 1B 02 AC 8A 21 01 30 00 00 00 02 
28 A3 02 2D 05 2A 02 A2 8C 01 28 C3 02 3D 05 3C 
02 C3 0E 49 C0 19 0C 2A 00 00 00 80 0E 24 C0 14 
98 01 9A 04 9C 04 0E 89 DB F5 01 20 00 00 00 00 
0E 29 C4 7D 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 0A 5C 0C 2D 00 00 00 04 92 01 
0E 28 C0 50 0B C9 0E 59 C3 E4 0C ED 00 00 00 04 
01 20 00 00 00 01 28 28 0C 3D 00 00 01 88 02 72 
26 73 0E 79 C0 29 0C 3D 00 00 01 8C 26 23 0E 29 
C4 3F 0C 20 00 00 00 0C 0A 3A 0D 04 FF FF FF DC 
0D 06 FF FF FF E0 0D 0E FF FF FF D8 19 50 0C 40 
FF FF FF DC 0C 60 FF FF FF E0 0C E0 FF FF FF D8 
0C 2D 00 00 00 04 0E 2E C7 8D 0A 26 0E 2D C3 B1 
1A 00 00 00 15 B2 0D 04 FF FF FF DC 0D 06 FF FF 
FF E0 0D 0E FF FF FF D8 19 50 0C 40 FF FF FF DC 
0C 60 FF FF FF E0 0C E0 FF FF FF D8 1A 00 00 00 
16 90 0D D8 00 00 00 04 1A 00 00 00 16 36 0A 2A 
0D 04 FF FF FF DC 0D 06 FF FF FF E0 0D 0E FF FF 
FF D8 19 50 0C E0 FF FF FF D8 0C 60 FF FF FF E0 
0C 40 FF FF FF DC 1A 00 00 00 16 90 0C 2D 00 00 
00 04 0E 29 C4 1B 0A 2D 0E 29 C0 1E 0B 62 02 2D 
0D 04 FF FF FF DC 0D 06 FF FF FF E0 03 00 00 00 
00 00 0C 60 FF FF FF E0 0A D6 0C 40 FF FF FF DC 
0E D9 C7 43 1A 00 00 00 16 14 0A 2D 02 6D 02 D2 
1A 00 00 00 17 40 02 29 1A 00 00 00 17 4C 06 18 
06 19 06 1A 06 1B 06 1C 06 1D 91 30 0D 02 00 00 
00 0C 02 83 0D 04 00 00 00 14 0C D4 00 00 00 08 
01 30 00 00 00 00 0E D3 C0 4A 38 28 00 00 00 0C 
01 50 00 00 00 10 02 42 28 45 27 45 01 50 00 00 
00 08 02 64 26 65 0E 63 C0 44 0C 58 00 00 00 10 
0E 53 C0 3F 0C 50 00 00 00 14 0A 95 01 50 00 00 
00 02 02 64 26 65 01 A0 00 00 00 00 0E 6A C0 57 
02 CA 02 DA 0E AD C0 AC 0C 38 00 00 00 1C 02 5A 
01 70 00 00 04 00 0E A7 E4 02 02 57 0C 68 00 00 
00 24 0C 20 00 00 00 0C 02 4C 19 60 0E 2D DC A7 
05 C2 29 A2 0C 40 00 00 00 14 0C 34 00 00 00 08 
29 32 0D 43 00 00 00 08 0E 3D C7 DD 02 2D 02 70 
97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 
0C 20 00 00 00 0C 02 38 03 00 00 00 31 F8 01 30 
00 00 00 00 0E 23 C0 04 1A 00 00 00 1D 72 38 28 
00 00 00 0C 01 30 00 00 00 10 02 42 28 43 27 43 
0C 50 00 00 00 14 0A 95 01 50 00 00 00 02 02 64 
26 65 01 A0 00 00 00 00 0E 6A C7 AB 01 30 00 00 
00 01 26 43 0E 46 C4 79 02 A4 02 D4 02 C4 0E AD 
C0 47 0C 58 00 00 00 08 01 60 00 00 00 10 28 26 
27 26 02 32 01 70 00 00 02 00 26 37 0E 3D C0 F9 
02 65 0E A5 E1 4D 02 BA 0A 28 02 6A 02 5A 02 3C 
02 46 0D 05 FF FF FF D8 0D 06 FF FF FF D0 01 70 
00 00 29 F8 19 70 0C 28 00 00 00 08 29 2B 0D 82 
00 00 00 08 0A 28 0C 60 FF FF FF D0 05 26 0B 82 
02 6A 0C 50 FF FF FF D8 05 C6 29 A6 0C 30 00 00 
00 14 0C 23 00 00 00 08 29 25 0D 32 00 00 00 08 
0E 2D C3 85 38 28 00 00 00 0C 0E AD C7 BB 0A C9 
0C A9 00 00 00 04 89 08 1A 00 00 00 18 8E 0A C9 
0C A9 00 00 00 04 89 08 1A 00 00 00 17 D4 01 20 
00 00 00 0C 0C 50 00 00 00 0C 0B 52 01 20 00 00 
00 40 38 58 00 00 00 0C 2B 25 39 82 00 00 00 0C 
01 20 FF FF FF FF 02 70 97 18 07 7D 07 7C 07 7B 
07 7A 07 79 07 78 04 00 0D 06 FF FF FF E0 02 C6 
02 D6 0D 06 FF FF FF E4 02 E6 0E CE C0 79 0C 60 
FF FF FF E0 0E 6E C0 4F 02 5D 0E DC E4 02 02 5C 
0C A8 00 00 00 08 0C 78 00 00 00 14 0D 07 FF FF 
FF DC 0A 28 0C 38 00 00 00 10 0E 23 E4 05 05 7A 
02 A7 0E 57 CD 5E 0C 70 FF FF FF DC 0E 57 C8 88 
0C 68 00 00 00 24 0C 20 00 00 00 0C 0C 38 00 00 
00 1C 0C 40 FF FF FF E4 02 57 0D 0E FF FF FF D4 
19 60 02 A2 0C E0 FF FF FF D4 0E 2E DF A8 29 DA 
0E DE C0 90 0C 30 FF FF FF E4 05 3A 0D 03 FF FF 
FF E4 29 CA 0C 40 00 00 00 14 0C 24 00 00 00 08 
29 2A 0D 42 00 00 00 08 0E 2E C7 B0 02 2E 1A 00 
00 00 18 1E 0C 20 FF FF FF E4 01 30 00 00 00 0A 
02 4C 0D 0E FF FF FF D4 01 70 00 00 27 E4 19 70 
0C 30 FF FF FF E0 0E 23 0C E0 FF FF FF D4 C1 7F 
02 D2 8D 01 0C 40 FF FF FF E4 29 D4 01 50 00 00 
00 01 0D 05 FF FF FF E0 1A 00 00 00 19 98 0A 49 
0D 04 FF FF FF E4 0C C9 00 00 00 04 89 08 01 50 
00 00 00 00 0D 05 FF FF FF E0 1A 00 00 00 19 8A 
0A 28 0C 38 00 00 00 10 0E 23 E4 03 0E A5 D5 07 
0C 58 00 00 00 14 0E A5 D0 58 0C 68 00 00 00 24 
0C 20 00 00 00 0C 0C 38 00 00 00 1C 02 4C 19 60 
02 52 0E 2D DF 3C 02 62 1A 00 00 00 18 F8 0C 30 
FF FF FF E4 02 45 0D 05 FF FF FF D8 0D 0E FF FF 
FF D4 01 60 00 00 29 F8 19 60 0C 28 00 00 00 08 
0C 50 FF FF FF D8 29 25 0D 82 00 00 00 08 0A 28 
05 25 0B 82 02 A5 0C E0 FF FF FF D4 29 DA 0E DE 
C7 72 0C 20 00 00 00 0C 02 38 0D 0E FF FF FF D4 
01 70 00 00 33 C0 19 70 0E 2D 0C E0 FF FF FF D4 
C7 06 0D 0D FF FF FF E0 1A 00 00 00 1A 04 02 32 
01 40 00 00 04 80 26 34 0E 3D C4 21 0A 28 02 B5 
02 5A 1A 00 00 00 18 BE 02 3C 02 4A 0D 0A FF FF 
FF D8 01 60 00 00 29 F8 19 60 0C 28 00 00 00 08 
29 2A 0D 82 00 00 00 08 0A 28 05 2A 0B 82 02 6A 
0C 50 FF FF FF D8 1A 00 00 00 18 F8 0C 38 00 00 
00 10 0A 68 29 63 0C 58 00 00 00 14 02 45 05 45 
05 45 02 54 01 70 00 00 00 1F 27 57 05 54 01 40 
00 00 00 01 2D 54 02 45 02 76 87 01 05 7A 0E 57 
E0 03 02 57 02 47 01 70 00 00 04 00 26 27 0E 2D 
C0 96 0C 20 00 00 00 0C 02 34 0D 05 FF FF FF D8 
0D 06 FF FF FF D0 03 00 00 00 1D A0 0E 2D 0C 50 
FF FF FF D8 0C 60 FF FF FF D0 C2 9A 0C 38 00 00 
00 10 02 46 0D 05 FF FF FF D8 0D 06 FF FF FF D0 
0D 02 FF FF FF D4 03 00 00 00 29 06 01 20 FF FF 
FB 7F 38 78 00 00 00 0C 26 27 01 30 00 00 00 80 
2B 23 39 82 00 00 00 0C 0C 50 FF FF FF D8 0C 60 
FF FF FF D0 0C E0 FF FF FF D4 0D 8E 00 00 00 10 
02 2E 05 26 0B 82 0D 85 00 00 00 14 02 BA 29 56 
0D 85 00 00 00 08 02 6A 02 5A 1A 00 00 00 18 BE 
0C 30 FF FF FF E4 02 47 0D 0E FF FF FF D4 01 50 
00 00 29 F8 19 50 0A 28 05 2A 0B 82 0C 20 00 00 
00 0C 02 38 01 60 00 00 33 C0 19 60 0C E0 FF FF 
FF D4 0E 2E C2 A5 1A 00 00 00 19 4C 02 3C 02 45 
0D 05 FF FF FF D8 0D 05 FF FF FF D0 01 70 00 00 
29 F8 19 70 0A 28 0C 50 FF FF FF D8 05 25 0B 82 
0C 20 00 00 00 0C 02 38 01 40 00 00 33 C0 19 40 
0E 2D 0C 50 FF FF FF D8 0C 60 FF FF FF D0 C4 04 
1A 00 00 00 18 F8 1A 00 00 00 19 4C 0C 20 00 00 
00 0C 0D 05 FF FF FF D8 0D 06 FF FF FF D0 03 00 
00 00 2B 36 02 E2 0E 2D 0C 50 FF FF FF D8 0C 60 
FF FF FF D0 C7 93 0C 20 00 00 00 0C 0C 38 00 00 
00 10 03 00 00 00 3B A0 01 20 00 00 00 0C 0C 30 
00 00 00 0C 0B 32 1A 00 00 00 19 4C 02 DC 8D 01 
01 60 00 00 00 01 0D 06 FF FF FF E0 1A 00 00 00 
19 98 01 20 00 00 00 40 38 38 00 00 00 0C 2B 23 
39 82 00 00 00 0C 01 20 00 00 00 09 0C 40 00 00 
00 0C 0B 42 01 20 FF FF FF FF 1A 00 00 00 18 1E 
06 18 06 19 06 1A 06 1B 06 1C 06 1D 91 28 02 92 
02 83 88 0B 01 20 00 00 00 16 0E 82 E4 59 01 20 
FF FF FF F8 26 82 01 20 00 00 00 00 0E 82 C8 55 
0E 38 D4 53 02 29 03 00 00 00 2B 32 01 20 00 00 
01 F7 0E 82 D4 5A 01 20 00 00 00 03 02 68 27 62 
01 30 00 00 4F 5C 0D 03 FF FF FF E4 02 46 28 42 
05 34 0C A3 00 00 00 0C 0E A3 C4 04 1A 00 00 00 
24 E4 0C 2A 00 00 00 04 01 30 FF FF FF FC 26 23 
0C 3A 00 00 00 0C 0C 4A 00 00 00 08 0D 43 00 00 
00 0C 0D 34 00 00 00 08 02 3A 05 32 0C 23 00 00 
00 04 01 40 00 00 00 01 2B 24 0D 32 00 00 00 04 
02 29 03 00 00 00 2B 34 02 2A 82 08 02 70 97 18 
07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 01 80 
00 00 00 10 0E 38 E7 AF 01 20 00 00 00 0C 0B 92 
01 20 00 00 00 00 02 70 97 18 07 7D 07 7C 07 7B 
07 7A 07 79 07 78 04 00 01 60 00 00 00 09 02 58 
27 56 02 65 01 20 00 00 00 00 0E 52 C1 36 01 20 
00 00 00 04 0E 52 E4 04 1A 00 00 00 24 7E 01 60 
00 00 00 06 02 28 27 26 02 62 86 38 01 40 00 00 
00 03 02 36 28 34 02 43 01 30 00 00 4F 5C 0D 03 
FF FF FF E4 05 34 02 43 0C A3 00 00 00 0C 0E 3A 
C0 2F 0C 2A 00 00 00 04 01 70 FF FF FF FC 26 27 
02 32 29 38 01 50 00 00 00 0F 0E 35 DC 04 1A 00 
00 00 23 D4 01 C0 00 00 00 00 0E 3C C8 14 1A 00 
00 00 23 DC 0C 2A 00 00 00 04 26 27 02 32 29 38 
0E 35 DC 04 1A 00 00 00 23 D4 0E 3C C8 04 1A 00 
00 00 23 DC 0C AA 00 00 00 0C 0E 4A C7 EC 86 01 
01 40 00 00 4F 64 08 A0 00 00 4F 6C 0E 4A C1 39 
0C 2A 00 00 00 04 01 30 FF FF FF FC 26 23 02 32 
29 38 01 50 00 00 00 0F 0E 35 DC 04 1A 00 00 00 
24 B2 0D 44 00 00 00 0C 0D 44 00 00 00 08 01 70 
00 00 00 00 0E 37 C8 04 1A 00 00 00 24 2C 01 30 
00 00 01 FF 0E 23 D4 C4 01 50 00 00 00 03 27 25 
01 70 00 00 00 02 02 32 2D 37 02 73 01 30 00 00 
00 01 28 37 08 70 00 00 4F 60 2B 37 0C 70 FF FF 
FF E4 0D 73 00 00 00 04 28 25 05 72 0C 57 00 00 
00 08 0D A7 00 00 00 0C 0D A5 00 00 00 08 0D 7A 
00 00 00 08 0D 5A 00 00 00 0C 01 20 00 00 00 02 
02 76 2D 72 01 50 00 00 00 01 28 57 0E 53 D4 EF 
02 73 26 75 01 20 00 00 00 00 0E 72 C4 11 01 20 
FF FF FF FC 26 62 86 04 05 55 02 23 26 25 0E 27 
C4 07 86 04 05 55 02 75 26 73 0E 72 C3 FB 01 C0 
FF FF FF FC 01 D0 00 00 00 0F 01 E0 00 00 00 00 
0D 05 FF FF FF DC 02 26 01 30 00 00 00 03 28 23 
0C 50 FF FF FF E4 05 52 0D 05 FF FF FF E0 02 76 
0C A5 00 00 00 0C 0E 5A C4 11 1A 00 00 00 24 CA 
0E 3E C8 04 1A 00 00 00 25 00 0C AA 00 00 00 0C 
0E 5A C4 04 1A 00 00 00 24 CA 0C 2A 00 00 00 04 
26 2C 02 32 29 38 0E 3D DF EC 02 2A 05 28 01 50 
00 00 00 01 2B 85 0D A8 00 00 00 04 0C 6A 00 00 
00 0C 0C 8A 00 00 00 08 0D 86 00 00 00 0C 0D 68 
00 00 00 08 0D 42 00 00 00 0C 0D 42 00 00 00 08 
0D 24 00 00 00 0C 0D 24 00 00 00 08 02 63 2B 65 
0D 26 00 00 00 04 05 23 0B 23 02 29 03 00 00 00 
2B 34 02 2A 82 08 02 70 97 18 07 7D 07 7C 07 7B 
07 7A 07 79 07 78 04 00 01 40 00 00 00 03 02 68 
27 64 02 76 28 74 02 47 1A 00 00 00 1E D8 01 30 
00 00 00 09 02 72 27 73 02 37 01 70 00 00 00 04 
0E 37 D4 04 1A 00 00 00 25 56 01 70 00 00 00 14 
0E 37 E4 04 1A 00 00 00 26 58 02 73 87 5B 01 50 
00 00 00 03 02 37 28 35 02 53 0C 30 FF FF FF E4 
05 35 02 53 0C 33 00 00 00 08 0E 35 C4 04 1A 00 
00 00 25 E8 0C C3 00 00 00 04 01 70 FF FF FF FC 
26 C7 0E 2C D0 0A 1A 00 00 00 21 B2 0C C3 00 00 
00 04 26 C7 0E 2C E0 06 0C 33 00 00 00 08 0E 53 
C7 F6 0C 23 00 00 00 0C 0D A2 00 00 00 0C 0D A3 
00 00 00 08 0D 2A 00 00 00 08 0D 3A 00 00 00 0C 
08 30 00 00 4F 60 01 20 00 00 00 02 02 76 2D 72 
01 50 00 00 00 01 28 57 0E 53 E7 13 08 A0 00 00 
4F 64 0C DA 00 00 00 04 01 20 FF FF FF FC 26 D2 
0E 8D D4 08 02 2D 29 28 01 30 00 00 00 0F 0E 23 
CD 14 08 C0 00 00 53 8C 8C 10 05 C8 01 20 FF FF 
FF FF 08 30 00 00 53 68 0E 32 C0 09 01 20 00 00 
0F FF 05 C2 01 20 FF FF F0 00 26 C2 01 50 00 00 
31 AC 02 29 02 3C 0D 05 FF FF FF D8 19 50 02 42 
01 30 FF FF FF FF 0E 23 0C 50 FF FF FF D8 C1 91 
02 6A 05 6D 0E 62 D5 88 08 30 00 00 53 98 02 7C 
05 73 02 37 09 70 00 00 53 98 0E 62 C4 04 1A 00 
00 00 26 FC 01 70 FF FF FF FF 08 E0 00 00 53 68 
0E E7 C4 04 1A 00 00 00 27 46 02 72 05 73 02 37 
29 36 09 30 00 00 53 98 01 30 00 00 00 07 02 62 
26 63 02 36 01 60 00 00 00 00 0E 36 C1 90 01 60 
00 00 00 08 29 63 02 42 05 46 01 20 00 00 10 00 
05 62 02 24 05 2C 01 30 00 00 0F FF 26 23 02 C6 
29 C2 02 29 02 3C 0D 04 FF FF FF D8 19 50 01 30 
FF FF FF FF 0E 23 0C 40 FF FF FF D8 C4 04 1A 00 
00 00 27 52 29 24 05 2C 01 30 00 00 00 01 2B 23 
08 30 00 00 53 98 05 C3 02 3C 09 C0 00 00 53 98 
0C 70 FF FF FF E4 0D 74 00 00 00 08 0D 42 00 00 
00 04 0E 7A C0 24 01 20 00 00 00 0F 0E D2 E5 6B 
9D 0C 01 40 FF FF FF F8 26 D4 02 4A 05 4D 01 50 
00 00 00 05 0D 45 00 00 00 04 0D 45 00 00 00 08 
0C 4A 00 00 00 04 01 50 00 00 00 01 26 45 02 5D 
2B 54 0D A5 00 00 00 04 0E D2 D5 10 08 A0 00 00 
4F 64 08 20 00 00 53 90 0E 32 E4 04 09 30 00 00 
53 90 08 20 00 00 53 94 0E 32 E4 04 09 30 00 00 
53 94 0C 2A 00 00 00 04 01 30 FF FF FF FC 26 23 
0E 82 D4 07 29 28 01 30 00 00 00 0F 0E 23 CC 3D 
02 29 03 00 00 00 2B 34 01 20 00 00 00 00 1A 00 
00 00 1E 5C 96 01 1A 00 00 00 1F 4E 0C 3A 00 00 
00 0C 0C 4A 00 00 00 08 0D 43 00 00 00 0C 0D 34 
00 00 00 08 02 4A 05 42 02 24 0C 32 00 00 00 04 
01 40 00 00 00 01 2B 34 0D 23 00 00 00 04 02 29 
03 00 00 00 2B 34 02 2A 82 08 02 70 97 18 07 7D 
07 7C 07 7B 07 7A 07 79 07 78 04 00 02 7A 05 72 
02 27 1A 00 00 00 23 FA 01 30 00 00 00 01 02 48 
2B 43 0D A4 00 00 00 04 02 6A 05 68 0C 70 FF FF 
FF E4 0D 76 00 00 00 08 2B 23 0D 62 00 00 00 04 
02 29 03 00 00 00 2B 34 02 2A 82 08 02 70 97 18 
07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 01 20 
00 00 00 14 0E 52 E4 5E 01 20 00 00 00 54 0E 52 
D4 91 01 60 00 00 00 0C 02 78 27 76 02 67 86 6E 
01 40 00 00 00 03 02 26 28 24 02 42 1A 00 00 00 
1E D8 02 2A 05 28 01 50 00 00 00 01 2B 85 0D A8 
00 00 00 04 1A 00 00 00 20 D4 87 01 02 27 01 30 
00 00 00 03 26 23 0E 2E C0 D5 02 5A 85 08 1A 00 
00 00 20 70 02 2A 82 08 0C A2 00 00 00 0C 0E 2A 
C0 04 1A 00 00 00 1E 12 86 02 1A 00 00 00 1F 50 
02 7A 05 72 0C 37 00 00 00 04 01 40 00 00 00 01 
2B 34 0D 73 00 00 00 04 0C 2A 00 00 00 0C 0C 3A 
00 00 00 08 0D 32 00 00 00 0C 0D 23 00 00 00 08 
02 29 03 00 00 00 2B 34 02 2A 82 08 1A 00 00 00 
1E 5C 86 5B 01 40 00 00 00 03 02 56 28 54 02 45 
1A 00 00 00 1E D8 01 70 00 00 00 06 02 32 27 37 
02 73 87 38 01 50 00 00 00 03 02 37 28 35 02 53 
1A 00 00 00 21 6A 0C 70 FF FF FF E4 0E 7A C2 75 
08 A0 00 00 4F 64 0C 2A 00 00 00 04 01 30 FF FF 
FF FC 26 23 1A 00 00 00 23 B0 02 29 02 3A 83 08 
03 00 00 00 3B A0 08 30 00 00 53 98 1A 00 00 00 
23 7C 01 20 00 00 01 54 0E 52 D4 3A 01 60 00 00 
00 0F 02 38 27 36 02 63 86 77 01 40 00 00 00 03 
02 56 28 54 02 45 1A 00 00 00 1E D8 01 60 00 00 
10 00 1A 00 00 00 22 D2 01 20 00 00 00 02 2D 72 
01 C0 00 00 00 01 28 C7 08 20 00 00 4F 60 2B 2C 
0C 50 FF FF FF E4 0D 52 00 00 00 04 02 23 1A 00 
00 00 21 B8 01 20 00 00 00 01 0D 42 00 00 00 04 
02 A4 01 20 00 00 00 00 1A 00 00 00 23 B0 01 20 
00 00 05 54 0E 52 D4 7F 01 60 00 00 00 12 02 78 
27 76 02 67 86 7C 01 40 00 00 00 03 02 26 28 24 
02 42 1A 00 00 00 1E D8 01 70 00 00 00 54 0E 37 
D4 82 01 70 00 00 00 0C 02 52 27 57 02 75 87 6E 
01 50 00 00 00 03 02 37 28 35 02 53 1A 00 00 00 
21 6A 0C 20 FF FF FF E0 1A 00 00 00 26 90 96 01 
02 36 01 50 00 00 00 03 26 35 0E 3E C0 8A 02 32 
93 08 0A 22 0E 23 C3 F4 08 20 00 00 4F 60 0C 50 
FF FF FF DC 05 55 0D 05 FF FF FF DC 0E 52 E4 04 
1A 00 00 00 21 EC 0E 5E C4 04 1A 00 00 00 21 EC 
02 32 26 35 0E 3E C0 05 02 67 1A 00 00 00 20 56 
02 35 87 04 05 33 02 53 26 52 0E 5E C3 FB 0D 03 
FF FF FF DC 02 67 1A 00 00 00 20 56 01 E0 00 00 
0F FF 02 76 26 7E 02 E7 01 70 00 00 00 00 0E E7 
C0 04 1A 00 00 00 22 84 08 A0 00 00 4F 64 05 CD 
01 20 00 00 00 01 2B C2 0D AC 00 00 00 04 1A 00 
00 00 23 82 01 40 00 00 03 F0 01 60 00 00 00 7E 
1A 00 00 00 1E D8 09 20 00 00 53 68 1A 00 00 00 
22 A8 01 20 00 00 00 01 01 C0 00 00 00 00 1A 00 
00 00 23 10 01 70 00 00 01 54 0E 37 D4 0D 02 72 
27 75 87 77 01 50 00 00 00 03 02 37 28 35 02 53 
1A 00 00 00 21 6A 01 50 00 00 05 54 0E 35 D4 22 
01 70 00 00 00 12 02 52 27 57 02 75 87 7C 01 50 
00 00 00 03 02 37 28 35 02 53 1A 00 00 00 21 6A 
0C 60 FF FF FF DC 2C 26 08 30 00 00 4F 60 26 23 
0C 30 FF FF FF E4 0D 32 00 00 00 04 1A 00 00 00 
26 AE 01 50 00 00 03 F0 01 70 00 00 00 7E 1A 00 
00 00 21 6A 06 18 06 19 06 1A 06 1B 06 1C 02 52 
02 93 01 80 00 00 00 03 02 A2 26 A8 01 60 00 00 
00 00 0E A6 C0 23 0E 46 C0 76 01 E0 00 00 00 18 
1C B2 28 BE 27 BE 02 A3 28 AE 27 AE 0E BA C0 63 
94 01 02 2E 02 E9 28 E2 27 E2 1A 00 00 00 28 40 
0E 46 C0 61 1C A5 28 A2 27 A2 0E AE C0 53 94 01 
85 01 02 A5 26 A8 0E A6 C7 F4 01 E0 00 00 00 03 
0E 4E E4 2C 01 60 00 00 00 18 02 23 28 26 27 26 
01 60 00 00 00 08 02 82 28 86 02 68 2B 62 01 20 
00 00 00 10 02 B6 28 B2 02 2B 2B 26 01 A0 FE FE 
FE FF 01 80 80 80 80 80 01 60 00 00 00 00 0A C5 
02 B2 2E BC 02 CB 05 BA 2C CC 26 BC 26 B8 0E B6 
C4 05 94 04 85 04 0E 4E D7 F3 01 60 00 00 00 00 
0E 46 C0 21 01 20 00 00 00 18 1C 85 28 82 27 82 
28 32 27 32 0E 83 C0 0E 94 01 02 36 28 92 27 92 
0E 43 C0 11 85 01 94 01 1C 65 28 62 27 62 0E 69 
C7 F8 02 25 02 70 97 14 07 7C 07 7B 07 7A 07 79 
07 78 04 00 02 24 02 70 97 14 07 7C 07 7B 07 7A 
07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 02 62 
02 E3 02 54 01 80 00 00 00 0F 0E 48 E4 59 02 93 
2B 92 01 A0 00 00 00 03 26 9A 01 A0 00 00 00 00 
0E 9A C4 4E 02 E4 02 63 02 52 0A 96 0B 59 0C 96 
00 00 00 04 0D 59 00 00 00 04 0C 96 00 00 00 08 
0D 59 00 00 00 08 0C 96 00 00 00 0C 0D 59 00 00 
00 0C 85 10 86 10 9E 10 0E E8 D7 E8 94 10 01 80 
00 00 00 04 02 54 27 58 02 E5 8E 01 28 E8 02 62 
05 6E 05 3E 02 E3 28 58 29 45 02 54 01 30 00 00 
00 03 0E 43 E4 1D 01 50 00 00 00 00 02 86 05 85 
02 9E 05 95 0A 99 0B 89 85 04 02 84 29 85 0E 83 
D7 F6 94 04 01 80 00 00 00 02 02 54 27 58 02 35 
83 01 28 38 05 63 05 E3 28 58 29 45 02 54 01 40 
00 00 00 00 0E 54 C0 0A 02 36 05 34 02 8E 05 84 
1C 88 1E 38 84 01 0E 45 C7 F8 02 70 97 10 07 7B 
07 7A 07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 
02 62 02 E3 02 54 0E 23 E4 1E 02 83 05 84 0E 28 
E0 1A 01 30 00 00 00 00 0E 43 C0 0E 02 32 05 34 
94 01 01 50 FF FF FF FF 93 01 98 01 1C 68 1E 36 
94 01 0E 45 C7 FA 02 70 97 10 07 7B 07 7A 07 79 
07 78 04 00 01 80 00 00 00 0F 0E 48 D4 16 01 40 
00 00 00 00 0E 54 C3 F0 02 36 05 34 02 8E 05 84 
1C 88 1E 38 84 01 0E 45 C7 F8 02 70 97 10 07 7B 
07 7A 07 79 07 78 04 00 02 93 2B 92 01 A0 00 00 
00 03 26 9A 01 A0 00 00 00 00 0E 9A C7 E1 02 E4 
02 63 02 52 0A 96 0B 59 0C 96 00 00 00 04 0D 59 
00 00 00 04 0C 96 00 00 00 08 0D 59 00 00 00 08 
0C 96 00 00 00 0C 0D 59 00 00 00 0C 85 10 86 10 
9E 10 0E E8 D7 E8 94 10 01 80 00 00 00 04 02 54 
27 58 02 E5 8E 01 28 E8 02 62 05 6E 05 3E 02 E3 
28 58 02 34 29 35 02 53 01 80 00 00 00 03 0E 38 
E7 AF 01 40 00 00 00 00 02 58 02 86 05 84 02 9E 
05 94 0A 99 0B 89 84 04 02 83 29 84 0E 85 D7 F6 
93 04 01 90 00 00 00 02 02 53 27 59 02 85 88 01 
28 89 05 68 05 E8 28 59 29 35 02 53 1A 00 00 00 
2A 4E 04 00 04 00 06 18 06 19 06 1A 06 1B 06 1C 
06 1D 91 24 0D 02 00 00 00 0C 02 93 01 A0 00 00 
00 00 0E 3A C1 C8 0D 04 FF FF FF E0 03 00 00 00 
2B 32 02 C9 9C 08 0C 5C 00 00 00 04 0C 40 FF FF 
FF E0 02 84 88 0B 01 20 00 00 00 16 0E 82 E4 BD 
01 20 FF FF FF F8 26 82 02 28 0E 8A C8 FF 0E 48 
D4 FD 01 70 FF FF FF FC 02 D5 26 D7 0E D2 D8 B4 
02 3C 05 3D 08 B0 00 00 4F 64 0D 0B FF FF FF E4 
0E B3 C1 A8 0C A3 00 00 00 04 01 60 FF FF FF FE 
02 BA 26 B6 02 6B 02 B3 05 B6 0C EB 00 00 00 04 
01 60 00 00 00 01 26 E6 01 60 00 00 00 00 0E E6 
C0 BE 02 36 01 70 00 00 00 01 26 57 02 75 01 50 
00 00 00 00 0E 75 C5 04 0A EC 02 5C 29 5E 02 E5 
0C 55 00 00 00 04 01 A0 FF FF FF FC 26 5A 0E 37 
C0 F3 0C 70 FF FF FF E4 0E 37 C4 04 1A 00 00 00 
30 24 02 75 05 7D 02 A6 05 A7 0E A2 C8 E7 0C 23 
00 00 00 0C 0C 33 00 00 00 08 0D 32 00 00 00 0C 
0D 23 00 00 00 08 0C 2E 00 00 00 0C 0C 3E 00 00 
00 08 0D 32 00 00 00 0C 0D 23 00 00 00 08 02 CE 
8C 08 9D 04 01 30 00 00 00 24 0E D3 E4 04 1A 00 
00 00 31 24 02 2C 01 40 00 00 00 13 0E D4 E4 29 
0A 29 0B C2 0C 29 00 00 00 04 0D E2 00 00 00 0C 
02 2E 82 10 89 08 01 40 00 00 00 1B 0E D4 E4 19 
0A 49 0B 24 0C 29 00 00 00 04 0D E2 00 00 00 14 
02 2E 82 18 89 08 0E D3 C4 0C 0A 39 0B 23 0C 29 
00 00 00 04 0D E2 00 00 00 1C 02 2E 82 20 89 08 
0A 39 0B 23 82 04 89 04 0A 39 0B 23 0C 39 00 00 
00 04 0D 23 00 00 00 04 0C 5E 00 00 00 04 02 9C 
02 CE 1A 00 00 00 2D 0C 01 20 00 00 00 10 02 82 
1A 00 00 00 2B 8E 02 9C 89 08 02 AD 02 2A 29 28 
01 30 00 00 00 0F 0E 23 D4 4D 01 30 00 00 00 01 
26 53 2B 5A 0D C5 00 00 00 04 05 CA 0C 2C 00 00 
00 04 2B 23 0D C2 00 00 00 04 0C 20 00 00 00 0C 
03 00 00 00 2B 34 02 A9 02 2A 02 70 97 18 07 7D 
07 7C 07 7B 07 7A 07 79 07 78 04 00 02 6A 26 67 
02 A6 05 AD 0E A2 CB 3F 0C 23 00 00 00 0C 0C 33 
00 00 00 08 0D 32 00 00 00 0C 0D 23 00 00 00 08 
02 9C 89 08 1A 00 00 00 2D 0C 01 20 00 00 00 0C 
0C 60 00 00 00 0C 0B 62 01 A0 00 00 00 00 02 2A 
02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 
04 00 02 3C 05 38 01 60 00 00 00 01 26 56 2B 58 
0D C5 00 00 00 04 02 42 2B 46 0D 34 00 00 00 04 
02 73 05 72 0C 47 00 00 00 04 2B 46 0D 74 00 00 
00 04 0C 20 00 00 00 0C 83 08 03 00 00 00 3B A0 
1A 00 00 00 2D 3A 02 75 05 7D 0E 72 D8 96 0C 20 
00 00 00 0C 02 34 03 00 00 00 1D A0 02 A2 01 30 
00 00 00 00 0E 23 C0 57 02 32 93 08 0C 5C 00 00 
00 04 01 40 FF FF FF FE 02 B5 26 B4 02 6C 05 6B 
0E 36 C1 6C 9D 04 01 30 00 00 00 24 0E D3 D4 EB 
02 29 02 4A 01 50 00 00 00 13 0E D5 E4 29 0A 29 
0B A2 0C 29 00 00 00 04 0D A2 00 00 00 04 84 08 
02 29 82 08 01 50 00 00 00 1B 0E D5 E4 19 0A 22 
0B 42 0C 29 00 00 00 0C 0D A2 00 00 00 0C 84 08 
02 29 82 10 0E D3 C4 0C 0A 22 0B 42 0C 29 00 00 
00 14 0D A2 00 00 00 14 84 08 02 29 82 18 0A 32 
0B 43 84 04 82 04 0A 32 0B 43 0C 22 00 00 00 04 
0D 42 00 00 00 04 0C 20 00 00 00 0C 02 39 03 00 
00 00 3B A0 0C 20 00 00 00 0C 03 00 00 00 2B 34 
02 2A 02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 
07 78 04 00 02 34 03 00 00 00 1D A0 02 A2 02 2A 
02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 
04 00 0C 30 FF FF FF E4 0C 63 00 00 00 04 26 67 
02 36 05 3D 02 78 87 10 0E 37 D8 5E 0C 30 FF FF 
FF E4 1A 00 00 00 2B E4 0C 2E 00 00 00 0C 0C 3E 
00 00 00 08 0D 32 00 00 00 0C 0D 23 00 00 00 08 
02 AE 8A 08 9D 04 01 30 00 00 00 24 0E D3 D4 FF 
02 2A 01 40 00 00 00 13 0E D4 E4 29 0A 29 0B A2 
0C 29 00 00 00 04 0D E2 00 00 00 0C 02 2E 82 10 
89 08 01 40 00 00 00 1B 0E D4 E4 19 0A 49 0B 24 
0C 29 00 00 00 04 0D E2 00 00 00 14 02 2E 82 18 
89 08 0E D3 C4 0C 0A 39 0B 23 0C 29 00 00 00 04 
0D E2 00 00 00 1C 02 2E 82 20 89 08 0A 39 0B 23 
82 04 89 04 0A 39 0B 23 0C 39 00 00 00 04 0D 23 
00 00 00 04 0C 5E 00 00 00 04 02 9A 02 A7 02 CE 
1A 00 00 00 2D 0C 02 2C 05 28 09 20 00 00 4F 64 
29 38 01 40 00 00 00 01 2B 34 0D 23 00 00 00 04 
0C 2C 00 00 00 04 26 24 2B 82 0D C8 00 00 00 04 
0C 20 00 00 00 0C 03 00 00 00 2B 34 02 A9 1A 00 
00 00 2D 48 02 39 02 4D 03 00 00 00 29 F8 1A 00 
00 00 2E B6 02 75 05 7D 05 67 02 38 83 10 0E 63 
CA E5 0C 2E 00 00 00 0C 0C 3E 00 00 00 08 0D 32 
00 00 00 0C 0D 23 00 00 00 08 02 AE 8A 08 9D 04 
01 30 00 00 00 24 0E D3 D4 95 02 2A 01 40 00 00 
00 13 0E D4 E4 29 0A 29 0B A2 0C 29 00 00 00 04 
0D E2 00 00 00 0C 02 2E 82 10 89 08 01 40 00 00 
00 1B 0E D4 E4 19 0A 49 0B 24 0C 29 00 00 00 04 
0D E2 00 00 00 14 02 2E 82 18 89 08 0E D3 C4 0C 
0A 39 0B 23 0C 29 00 00 00 04 0D E2 00 00 00 1C 
02 2E 82 20 89 08 0A 39 0B 23 82 04 89 04 0A 39 
0B 23 0C 39 00 00 00 04 0D 23 00 00 00 04 02 2E 
05 28 09 20 00 00 4F 64 29 68 01 30 00 00 00 01 
2B 63 0D 26 00 00 00 04 0C 2E 00 00 00 04 26 23 
2B 82 0D E8 00 00 00 04 0C 20 00 00 00 0C 03 00 
00 00 2B 34 1A 00 00 00 2D 48 0C A3 00 00 00 04 
01 20 FF FF FF FC 26 A2 05 AD 02 9C 89 08 1A 00 
00 00 2D 0C 02 2C 02 39 02 4D 0D 0E FF FF FF E0 
03 00 00 00 29 F8 0C E0 FF FF FF E0 0C 5E 00 00 
00 04 02 9C 02 CE 1A 00 00 00 2D 0C 02 2A 02 39 
02 4D 0D 07 FF FF FF DC 0D 0E FF FF FF E0 03 00 
00 00 29 F8 0C E0 FF FF FF E0 0C 5E 00 00 00 04 
02 9A 0C 70 FF FF FF DC 02 A7 02 CE 1A 00 00 00 
2D 0C 02 2A 02 39 02 4D 0D 06 FF FF FF DC 0D 0E 
FF FF FF E0 03 00 00 00 29 F8 0C E0 FF FF FF E0 
0C 60 FF FF FF DC 1A 00 00 00 30 CE 06 18 06 19 
06 1B 91 18 02 92 01 80 00 00 00 00 09 80 00 00 
53 C0 02 23 03 00 00 00 49 C4 01 30 FF FF FF FF 
0E 23 C0 07 02 70 97 0C 07 7B 07 79 07 78 04 00 
08 30 00 00 53 C0 0E 38 C3 F6 0B 93 02 70 97 0C 
07 7B 07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 
91 18 02 92 02 83 08 20 00 00 4B 34 01 30 00 00 
00 00 0E 23 C0 06 0C 42 00 00 00 38 0E 43 C0 68 
38 38 00 00 00 0C 02 E3 02 63 01 40 00 00 00 10 
02 23 28 24 27 24 01 50 00 00 00 08 02 A2 26 A5 
02 5A 01 A0 00 00 00 00 0E 5A C0 7B 0C 48 00 00 
00 10 01 20 00 00 00 00 0E 42 C0 50 01 20 00 00 
00 10 28 32 27 32 01 20 00 00 00 01 02 A3 26 A2 
02 2A 01 50 00 00 00 00 0E A5 C0 17 0D 85 00 00 
00 08 0C 28 00 00 00 14 2A 22 0D 82 00 00 00 18 
01 20 00 00 00 00 0E 42 C0 19 02 70 97 10 07 7B 
07 7A 07 79 07 78 04 00 01 50 00 00 00 02 26 35 
0E 3A C4 04 0C 28 00 00 00 14 0D 82 00 00 00 08 
01 20 00 00 00 00 0E 42 C7 E9 01 30 00 00 00 10 
38 28 00 00 00 0C 28 23 27 23 01 30 00 00 00 80 
26 23 0E 24 C4 28 02 24 1A 00 00 00 32 9A 03 00 
00 00 37 20 1A 00 00 00 32 20 01 50 00 00 00 10 
02 23 28 25 27 25 01 50 00 00 02 80 26 25 01 50 
00 00 02 00 0E 25 C3 A3 02 29 02 38 03 00 00 00 
40 AE 38 38 00 00 00 0C 0C 48 00 00 00 10 1A 00 
00 00 32 5C 01 20 FF FF FF FF 1A 00 00 00 32 9A 
02 32 26 34 0E 35 C3 F7 01 30 00 00 00 04 26 23 
0E 25 C4 10 0C 48 00 00 00 10 01 30 00 00 00 08 
02 56 2B 53 02 35 39 85 00 00 00 0C 1A 00 00 00 
32 52 0C 38 00 00 00 30 0E 35 C0 12 02 28 82 40 
0E 32 C0 08 02 29 03 00 00 00 3B A0 38 E8 00 00 
00 0C 01 20 00 00 00 00 0D 82 00 00 00 30 01 60 
FF FF FF DB 26 6E 01 20 00 00 00 00 0D 82 00 00 
00 04 0C 48 00 00 00 10 0B 84 1A 00 00 00 33 5A 
06 18 06 19 06 1A 06 1B 06 1C 06 1D 91 1C 02 C2 
02 83 01 30 00 00 00 00 0E 23 C0 06 0C 42 00 00 
00 38 0E 43 C0 E1 38 58 00 00 00 0C 01 20 00 00 
00 10 02 D5 28 D2 2D D2 01 40 00 00 00 00 0E D4 
C0 C9 01 A0 00 00 00 08 02 2D 26 2A 02 A2 0E 24 
C4 82 01 20 00 00 08 00 2B 52 39 85 00 00 00 0C 
0C 28 00 00 00 04 0E 2A DC F7 0C D8 00 00 00 28 
01 20 00 00 00 00 0E D2 C0 AD 01 90 00 00 00 10 
28 59 27 59 01 60 00 00 10 00 02 35 26 36 02 63 
0E 32 C0 B6 0C A8 00 00 00 50 01 20 00 00 00 04 
26 52 01 20 00 00 00 00 0E 52 C0 0E 0C 38 00 00 
00 04 29 A3 0C 38 00 00 00 30 0E 32 C0 05 0C 28 
00 00 00 3C 29 A2 02 2C 0C 38 00 00 00 1C 02 4A 
01 50 00 00 00 00 19 D0 0E A2 C4 66 01 20 FF FF 
F7 FF 38 38 00 00 00 0C 26 23 39 82 00 00 00 0C 
01 30 00 00 00 00 0D 83 00 00 00 04 0C 48 00 00 
00 10 0B 84 01 40 00 00 10 00 26 24 0E 23 C0 04 
0D 8A 00 00 00 50 0C 38 00 00 00 30 01 20 00 00 
00 00 0E 32 C0 A2 02 28 82 40 0E 32 C0 05 02 2C 
03 00 00 00 3B A0 01 20 00 00 00 00 0D 82 00 00 
00 30 02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 
07 78 04 00 0C A8 00 00 00 10 0E A4 C0 82 0A 98 
29 9A 0B 8A 01 20 00 00 00 03 26 D2 0E D4 C0 42 
0D 84 00 00 00 08 01 D0 00 00 00 00 0E 9D CC 08 
1A 00 00 00 35 92 29 92 0E 9D DC 5A 05 A2 0C 68 
00 00 00 24 02 2C 0C 38 00 00 00 1C 02 4A 02 59 
19 60 0E 2D CF F1 01 20 00 00 00 40 38 38 00 00 
00 0C 2B 23 39 82 00 00 00 0C 01 20 FF FF FF FF 
02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 
04 00 02 2D 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 03 00 00 00 37 20 1A 00 00 00 
33 E6 0C 48 00 00 00 14 1A 00 00 00 35 30 02 2C 
0C 38 00 00 00 1C 02 46 01 50 00 00 00 01 0D 06 
FF FF FF E4 19 D0 02 A2 01 20 FF FF FF FF 0E A2 
0C 60 FF FF FF E4 C0 25 38 58 00 00 00 0C 28 59 
27 59 0C D8 00 00 00 28 1A 00 00 00 34 5A 01 20 
00 00 00 00 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 0C 28 00 00 00 3C 0E 2A CF 06 
02 2A 1A 00 00 00 35 94 02 23 1A 00 00 00 35 94 
0A 3C 01 20 00 00 00 1D 0E 32 C0 0F 01 20 00 00 
00 40 38 38 00 00 00 0C 2B 23 39 82 00 00 00 0C 
02 2A 1A 00 00 00 35 94 02 26 1A 00 00 00 35 94 
06 1B 91 18 02 32 01 20 00 00 00 00 0E 32 C0 0B 
08 20 00 00 4B 34 03 00 00 00 33 C0 02 70 97 04 
07 7B 04 00 08 20 00 00 4A 24 01 30 00 00 33 C0 
03 00 00 00 3F CA 02 70 97 04 07 7B 04 00 01 20 
00 00 00 00 04 00 01 20 00 00 00 00 04 00 91 18 
01 30 00 00 48 1E 03 00 00 00 3E F8 04 00 06 18 
06 19 06 1A 06 1B 91 18 02 A3 01 90 00 00 00 68 
2F 39 02 93 83 0C 03 00 00 00 1D A0 02 82 01 30 
00 00 00 00 0E 23 C0 0D 82 0C 0B 83 0D 8A 00 00 
00 04 0D 82 00 00 00 08 02 49 03 00 00 00 11 6C 
02 28 02 70 97 10 07 7B 07 7A 07 79 07 78 04 00 
91 18 08 20 00 00 4A 24 03 00 00 00 36 AE 04 00 
06 18 06 19 06 1A 06 1B 06 1C 06 1D 91 20 02 92 
0C 82 00 00 00 38 01 20 00 00 00 00 0E 82 C4 E7 
01 20 00 00 36 AE 0D 92 00 00 00 3C 01 E0 00 00 
00 01 0D 9E 00 00 00 38 0D 98 00 00 02 E0 01 20 
00 00 00 03 0D 92 00 00 02 E4 01 20 00 00 02 EC 
02 39 05 32 0D 93 00 00 02 E8 0C A9 00 00 00 04 
0B A8 0D A8 00 00 00 04 0D A8 00 00 00 08 20 20 
00 00 00 04 39 A2 00 00 00 0C 0D A8 00 00 00 64 
39 A8 00 00 00 0E 0D A8 00 00 00 10 0D A8 00 00 
00 14 0D A8 00 00 00 18 01 C0 00 00 11 6C 02 2A 
82 5C 02 38 01 40 00 00 00 08 0D 0E FF FF FF E4 
19 C0 0D AA 00 00 00 1C 01 B0 00 00 44 B2 0D AB 
00 00 00 20 01 D0 00 00 45 18 0D AD 00 00 00 24 
01 50 00 00 45 A6 0D A5 00 00 00 28 01 60 00 00 
46 10 0D A6 00 00 00 2C 0C A9 00 00 00 08 0B A8 
0D A8 00 00 00 04 0D A8 00 00 00 08 20 20 00 00 
00 09 39 A2 00 00 00 0C 0D A8 00 00 00 64 0C E0 
FF FF FF E4 39 AE 00 00 00 0E 0D A8 00 00 00 10 
0D A8 00 00 00 14 0D A8 00 00 00 18 02 2A 82 5C 
02 38 01 40 00 00 00 08 0D 05 FF FF FF E4 0D 06 
FF FF FF E0 19 C0 0D AA 00 00 00 1C 0D AB 00 00 
00 20 0D AD 00 00 00 24 0C 50 FF FF FF E4 0D A5 
00 00 00 28 0C 60 FF FF FF E0 0D A6 00 00 00 2C 
0C 99 00 00 00 0C 0B 98 0D 98 00 00 00 04 0D 98 
00 00 00 08 20 20 00 00 00 12 39 92 00 00 00 0C 
0D 98 00 00 00 64 20 20 00 00 00 02 39 92 00 00 
00 0E 0D 98 00 00 00 10 0D 98 00 00 00 14 0D 98 
00 00 00 18 02 29 82 5C 02 38 01 40 00 00 00 08 
19 C0 0D 99 00 00 00 1C 0D 9B 00 00 00 20 0D 9D 
00 00 00 24 0C 50 FF FF FF E4 0D 95 00 00 00 28 
0C 60 FF FF FF E0 0D 96 00 00 00 2C 02 70 97 18 
07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 06 18 
06 19 06 1A 06 1B 06 1C 06 1D 91 1C 02 D2 08 C0 
00 00 4A 24 0C 3C 00 00 00 38 01 20 00 00 00 00 
0E 32 C0 6D 01 20 00 00 02 E0 05 C2 01 90 00 00 
00 00 01 A0 00 00 00 10 01 40 00 00 36 BE 0C 8C 
00 00 00 08 0C 2C 00 00 00 04 92 01 0E 29 D8 08 
1A 00 00 00 3A 0E 92 01 0E 29 C8 4A 88 68 38 38 
00 00 00 0C 28 3A 2D 3A 0E 39 C7 F6 20 20 FF FF 
FF FF 39 82 00 00 00 0E 20 20 00 00 00 01 39 82 
00 00 00 0C 01 90 00 00 00 00 0D 89 00 00 00 64 
0B 89 0D 89 00 00 00 08 0D 89 00 00 00 04 0D 89 
00 00 00 10 0D 89 00 00 00 14 0D 89 00 00 00 18 
02 28 82 5C 02 39 01 40 00 00 00 08 03 00 00 00 
11 6C 0D 89 00 00 00 30 0D 89 00 00 00 34 0D 89 
00 00 00 44 0D 89 00 00 00 48 02 28 02 70 97 18 
07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 0A 2C 
0E 29 C0 0C 02 C2 1A 00 00 00 39 5E 02 2C 03 00 
00 00 37 20 1A 00 00 00 39 44 02 2D 01 30 00 00 
00 04 0D 04 FF FF FF E4 19 40 0B C2 0E 29 0C 40 
FF FF FF E4 C7 E8 01 20 00 00 00 0C 0B D2 02 89 
1A 00 00 00 39 FA 04 00 04 00 04 00 04 00 91 18 
08 20 00 00 4B 34 01 30 00 00 36 9E 03 00 00 00 
3E F8 04 00 91 18 08 20 00 00 4B 34 01 30 00 00 
36 A6 03 00 00 00 3E F8 04 00 06 18 06 19 06 1A 
06 1B 06 1C 91 18 02 A2 02 C3 03 00 00 00 2B 32 
08 20 00 00 4F 64 0C 92 00 00 00 04 01 20 FF FF 
FF FC 26 92 01 80 00 00 0F EF 02 29 05 28 02 82 
29 8C 01 20 00 00 00 0C 27 82 98 01 28 82 01 20 
00 00 0F FF 0E 82 DC 0F 01 C0 00 00 31 AC 02 2A 
01 30 00 00 00 00 19 C0 08 30 00 00 4F 64 05 39 
0E 23 C0 10 02 2A 03 00 00 00 2B 34 01 20 00 00 
00 00 02 70 97 14 07 7C 07 7B 07 7A 07 79 07 78 
04 00 02 2A 2A 38 19 C0 01 30 FF FF FF FF 0E 23 
C0 20 29 98 01 C0 00 00 00 01 2B 9C 08 20 00 00 
4F 64 0D 29 00 00 00 04 08 20 00 00 53 98 29 28 
09 20 00 00 53 98 02 2A 03 00 00 00 2B 34 02 2C 
02 70 97 14 07 7C 07 7B 07 7A 07 79 07 78 04 00 
02 2A 01 30 00 00 00 00 19 C0 08 30 00 00 4F 64 
02 42 29 43 01 50 00 00 00 0F 0E 45 DF BC 08 50 
00 00 53 68 29 25 09 20 00 00 53 98 01 20 00 00 
00 01 2B 42 0D 34 00 00 00 04 1A 00 00 00 3A F4 
06 18 06 19 06 1A 06 1B 91 18 02 82 02 A3 01 90 
00 00 00 00 0E 39 C0 B8 03 00 00 00 2B 32 9A 08 
0C 5A 00 00 00 04 01 20 FF FF FF FE 02 35 26 32 
02 23 02 3A 05 32 0C 43 00 00 00 04 01 60 FF FF 
FF FC 26 46 01 60 00 00 4F 5C 08 70 00 00 4F 64 
0E 73 C0 E4 0D 34 00 00 00 04 01 70 00 00 00 01 
26 57 0E 59 C4 15 0A 9A 29 A9 05 29 0C 9A 00 00 
00 08 02 E6 8E 08 0E 9E C1 01 0C 7A 00 00 00 0C 
0D 97 00 00 00 0C 0D 79 00 00 00 08 02 95 02 53 
05 54 0C 55 00 00 00 04 01 70 00 00 00 01 26 57 
01 E0 00 00 00 00 0E 5E C4 10 05 24 0E 95 C0 73 
0C 43 00 00 00 08 0C 33 00 00 00 0C 0D 43 00 00 
00 0C 0D 34 00 00 00 08 01 30 00 00 00 01 02 42 
2B 43 0D A4 00 00 00 04 02 4A 05 42 0B 42 01 40 
00 00 00 00 0E 94 C4 4C 01 40 00 00 01 FF 0E 24 
E4 70 01 30 00 00 00 09 02 42 27 43 02 34 01 40 
00 00 00 04 0E 34 D4 BE 01 50 00 00 00 06 02 72 
27 75 02 57 85 38 01 40 00 00 00 03 02 35 28 34 
02 43 02 36 05 34 02 43 0C 33 00 00 00 08 0E 34 
C0 B9 0C 63 00 00 00 04 01 50 FF FF FF FC 26 65 
0E 26 D0 0A 1A 00 00 00 3D 00 0C 63 00 00 00 04 
26 65 0E 26 E0 06 0C 33 00 00 00 08 0E 43 C7 F6 
0C 23 00 00 00 0C 0D A2 00 00 00 0C 0D A3 00 00 
00 08 0D 2A 00 00 00 08 0D 3A 00 00 00 0C 02 28 
03 00 00 00 2B 34 02 70 97 10 07 7B 07 7A 07 79 
07 78 04 00 0C 43 00 00 00 08 01 50 00 00 4F 64 
0E 45 C7 8A 0D 4A 00 00 00 0C 0D 4A 00 00 00 08 
0D A4 00 00 00 0C 0D A4 00 00 00 08 02 32 2B 37 
0D A3 00 00 00 04 05 A2 0B A2 1A 00 00 00 3D 1E 
01 50 00 00 00 03 27 25 01 40 00 00 00 02 02 72 
2D 74 28 37 08 40 00 00 4F 60 2B 43 0D 64 00 00 
00 04 28 25 05 62 0C 26 00 00 00 08 0D A6 00 00 
00 0C 0D A2 00 00 00 08 0D 6A 00 00 00 08 0D 2A 
00 00 00 0C 1A 00 00 00 3D 1E 05 42 01 20 00 00 
00 01 26 52 0E 59 C4 10 0A 2A 29 A2 05 42 0C 2A 
00 00 00 0C 0C 3A 00 00 00 08 0D 32 00 00 00 0C 
0D 23 00 00 00 08 01 20 00 00 00 01 02 74 2B 72 
0D A7 00 00 00 04 0D 6A 00 00 00 08 08 20 00 00 
53 64 0E 42 D3 8D 02 28 08 30 00 00 53 8C 03 00 
00 00 3A 8A 1A 00 00 00 3D 1E 02 97 1A 00 00 00 
3C 2E 01 40 00 00 00 14 0E 34 D4 1F 02 53 85 5B 
01 40 00 00 00 03 02 75 28 74 02 47 1A 00 00 00 
3C C2 01 20 00 00 00 02 2D 52 01 40 00 00 00 01 
28 45 08 20 00 00 4F 60 2B 24 0D 62 00 00 00 04 
02 23 1A 00 00 00 3D 06 01 40 00 00 00 54 0E 34 
D4 11 01 50 00 00 00 0C 02 32 27 35 02 53 85 6E 
01 40 00 00 00 03 02 75 28 74 02 47 1A 00 00 00 
3C C2 01 40 00 00 01 54 0E 34 D4 11 01 50 00 00 
00 0F 02 32 27 35 02 53 85 77 01 40 00 00 00 03 
02 75 28 74 02 47 1A 00 00 00 3C C2 01 40 00 00 
05 54 0E 34 D4 11 01 50 00 00 00 12 02 32 27 35 
02 53 85 7C 01 40 00 00 00 03 02 75 28 74 02 47 
1A 00 00 00 3C C2 01 40 00 00 03 F0 01 50 00 00 
00 7E 1A 00 00 00 3C C2 06 18 06 19 06 1A 06 1B 
06 1C 06 1D 91 24 02 82 0D 03 00 00 00 10 03 00 
00 00 3A 56 01 20 00 00 02 E0 05 82 01 90 00 00 
00 00 0E 89 C0 4F 02 49 01 D0 00 00 00 10 01 60 
FF FF FF FF 0C 58 00 00 00 08 0C A8 00 00 00 04 
9A 01 0E A4 C8 2F 02 C5 8C 0C 1A 00 00 00 3F 52 
85 68 21 2C 28 2D 2D 2D 0E 24 C0 20 38 2C 00 00 
00 02 28 2D 2D 2D 0E 26 C0 19 02 25 0D 04 FF FF 
FF E0 0D 05 FF FF FF E4 0D 06 FF FF FF DC 0C 30 
00 00 00 10 19 30 2B 92 0C 60 FF FF FF DC 0C 50 
FF FF FF E4 0C 40 FF FF FF E0 9A 01 8C 68 0E A4 
DB D8 0A 88 0E 84 C7 C7 03 00 00 00 3A 58 02 29 
02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 
04 00 02 98 1A 00 00 00 3F A8 06 18 06 19 06 1A 
06 1B 06 1C 06 1D 91 24 0D 02 00 00 00 0C 0D 03 
00 00 00 10 03 00 00 00 3A 56 01 50 00 00 02 E0 
0C 20 00 00 00 0C 05 25 02 52 01 80 00 00 00 00 
0E 28 C0 52 02 D8 01 C0 00 00 00 10 01 60 FF FF 
FF FF 0C 45 00 00 00 08 0C 95 00 00 00 04 99 01 
0E 9D C8 32 02 A4 8A 0C 1A 00 00 00 40 30 84 68 
21 2A 28 2C 2D 2C 0E 2D C0 23 38 2A 00 00 00 02 
28 2C 2D 2C 0E 26 C0 1C 0C 20 00 00 00 0C 02 34 
0D 04 FF FF FF E0 0D 05 FF FF FF E4 0D 06 FF FF 
FF DC 0C 70 00 00 00 10 19 70 2B 82 0C 60 FF FF 
FF DC 0C 50 FF FF FF E4 0C 40 FF FF FF E0 99 01 
8A 68 0E 9D DB D5 0A 55 0E 5D C7 C4 03 00 00 00 
3A 58 02 28 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 02 82 1A 00 00 00 40 8C 06 18 
06 19 06 1A 06 1B 06 1C 06 1D 91 54 02 C2 02 83 
38 53 00 00 00 0C 01 90 00 00 00 10 02 45 28 49 
27 49 01 A0 00 00 00 02 02 34 26 3A 02 A3 01 30 
00 00 00 00 0E A3 C4 92 38 38 00 00 00 0E 28 39 
2D 39 0E 3A C8 5C 02 40 94 54 03 00 00 00 48 30 
0E 2A C8 4F 0C 20 FF FF FF B0 01 30 00 00 F0 00 
26 23 01 D0 00 00 00 01 01 30 00 00 20 00 0E 23 
C0 02 02 DA 01 30 00 00 80 00 0E 23 C0 AB 01 20 
00 00 08 00 38 38 00 00 00 0C 2B 23 39 82 00 00 
00 0C 01 A0 00 00 04 00 02 2C 02 3A 03 00 00 00 
1D A0 01 90 00 00 00 00 0E 29 C0 42 01 30 00 00 
36 AE 0D C3 00 00 00 3C 01 30 00 00 00 80 38 48 
00 00 00 0C 2B 34 39 83 00 00 00 0C 0B 82 0D 82 
00 00 00 10 0D 8A 00 00 00 14 0E D9 C4 54 02 70 
97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 
38 58 00 00 00 0C 02 45 28 49 27 49 01 20 00 00 
00 80 26 42 01 20 00 00 00 00 0E 42 C4 5D 01 A0 
00 00 04 00 01 20 00 00 08 00 2B 52 39 85 00 00 
00 0C 01 D0 00 00 00 00 1A 00 00 00 41 48 38 38 
00 00 00 0C 01 50 00 00 00 10 02 43 28 45 27 45 
01 50 00 00 02 00 26 45 0E 42 C7 CA 01 20 00 00 
00 02 2B 32 39 83 00 00 00 0C 02 28 82 43 0B 82 
0D 82 00 00 00 10 01 20 00 00 00 01 0D 82 00 00 
00 14 02 70 97 18 07 7D 07 7C 07 7B 07 7A 07 79 
07 78 04 00 01 40 00 00 00 10 38 38 00 00 00 0E 
28 34 02 2C 2D 34 03 00 00 00 48 7E 0E 29 C3 A0 
01 20 00 00 00 01 38 38 00 00 00 0C 2B 23 39 82 
00 00 00 0C 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 01 A0 00 00 00 40 1A 00 00 00 
41 C4 0C 38 00 00 00 28 01 20 00 00 45 A6 0E 32 
C7 4F 01 A0 00 00 04 00 02 2A 38 48 00 00 00 0C 
2B 24 39 82 00 00 00 0C 0D 8A 00 00 00 4C 1A 00 
00 00 41 48 06 18 06 19 06 1B 91 18 02 92 02 83 
0A 33 01 40 00 00 00 00 0E 34 C0 04 03 00 00 00 
42 B4 02 29 02 38 03 00 00 00 3B A0 02 70 97 0C 
07 7B 07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 
06 1C 06 1D 91 18 02 82 08 20 00 00 4B 34 0E 82 
C0 63 0C 48 00 00 00 4C 01 D0 00 00 00 00 0E 4D 
C0 1F 01 90 00 00 3B A0 02 CD 02 24 05 2D 0A 32 
0E 3C C4 05 1A 00 00 00 43 3C 02 3A 0A A3 02 28 
19 90 0E AC C7 FB 0C 48 00 00 00 4C 8D 04 01 20 
00 00 00 3C 0E D2 C7 EA 02 28 02 34 19 90 0C 38 
00 00 00 40 01 20 00 00 00 00 0E 32 C0 05 02 28 
03 00 00 00 3B A0 0C 38 00 00 01 48 01 20 00 00 
00 00 0E 32 C0 15 01 C0 00 00 01 4C 02 28 05 2C 
02 C2 0E 32 C0 0D 01 90 00 00 3B A0 1A 00 00 00 
43 94 02 3A 0A A3 02 28 19 90 0E CA C7 FB 0C 38 
00 00 00 54 01 20 00 00 00 00 0E 32 C0 05 02 28 
03 00 00 00 3B A0 0C 28 00 00 00 38 01 90 00 00 
00 00 0E 29 C4 0A 02 70 97 18 07 7D 07 7C 07 7B 
07 7A 07 79 07 78 04 00 0C 38 00 00 00 3C 02 28 
19 30 0C 38 00 00 02 E0 0E 39 C3 EE 02 28 03 00 
00 00 42 B4 02 70 97 18 07 7D 07 7C 07 7B 07 7A 
07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 06 1C 
06 1D 91 18 0D 02 00 00 00 0C 01 20 00 00 00 00 
0C 30 00 00 00 0C 0E 32 C0 3C 0C 30 00 00 00 0C 
0C C3 00 00 01 48 01 A0 00 00 00 00 0E CA C0 19 
01 D0 00 00 00 02 0C 9C 00 00 00 04 02 89 98 01 
0E 8A C8 0C 89 01 28 9D 02 2C 05 29 02 92 0A 29 
19 20 98 01 99 04 0E 8A DB FB 0A CC 0E CA C7 EC 
0C 20 00 00 00 0C 0C 32 00 00 00 3C 01 20 00 00 
00 00 0E 32 C0 05 0C 20 00 00 00 0C 19 30 02 70 
97 18 07 7D 07 7C 07 7B 07 7A 07 79 07 78 04 00 
08 20 00 00 4B 34 0D 02 00 00 00 0C 1A 00 00 00 
44 2A 06 18 06 1B 91 18 02 83 01 60 00 00 00 10 
38 33 00 00 00 0E 28 36 2D 36 03 00 00 00 49 1A 
01 30 00 00 00 00 0E 23 C8 0D 0C 38 00 00 00 50 
05 32 0D 83 00 00 00 50 02 70 97 08 07 7B 07 78 
04 00 01 30 FF FF EF FF 38 48 00 00 00 0C 26 34 
39 83 00 00 00 0C 02 70 97 08 07 7B 07 78 04 00 
01 20 00 00 00 00 04 00 06 18 06 19 06 1A 06 1B 
06 1C 91 18 02 C2 02 83 02 94 02 A5 38 53 00 00 
00 0C 01 60 00 00 00 10 02 35 28 36 27 36 01 40 
00 00 01 00 26 34 01 40 00 00 00 00 0E 34 C0 0F 
38 38 00 00 00 0E 28 36 2D 36 01 50 00 00 00 02 
03 00 00 00 48 CA 38 58 00 00 00 0C 01 20 FF FF 
EF FF 26 52 39 85 00 00 00 0C 01 40 00 00 00 10 
38 38 00 00 00 0E 28 34 02 2C 2D 34 02 49 02 5A 
03 00 00 00 46 2A 02 70 97 14 07 7C 07 7B 07 7A 
07 79 07 78 04 00 06 18 06 1B 91 18 02 83 01 60 
00 00 00 10 38 33 00 00 00 0E 28 36 2D 36 03 00 
00 00 48 CA 01 30 FF FF FF FF 0E 23 C0 13 01 30 
00 00 10 00 38 48 00 00 00 0C 2B 34 39 83 00 00 
00 0C 0D 82 00 00 00 50 02 70 97 08 07 7B 07 78 
04 00 01 30 FF FF EF FF 38 48 00 00 00 0C 26 34 
39 83 00 00 00 0C 02 70 97 08 07 7B 07 78 04 00 
91 18 01 40 00 00 00 10 38 33 00 00 00 0E 28 34 
2D 34 03 00 00 00 46 7A 04 00 06 18 06 19 06 1B 
91 18 02 92 01 80 00 00 00 00 09 80 00 00 53 C0 
02 23 02 34 02 45 03 00 00 00 49 F6 01 30 FF FF 
FF FF 0E 23 C0 07 02 70 97 0C 07 7B 07 79 07 78 
04 00 08 30 00 00 53 C0 0E 38 C3 F6 0B 93 02 70 
97 0C 07 7B 07 79 07 78 04 00 06 18 06 19 06 1B 
91 18 02 92 01 80 00 00 00 00 09 80 00 00 53 C0 
02 23 03 00 00 00 49 D8 01 30 FF FF FF FF 0E 23 
C0 07 02 70 97 0C 07 7B 07 79 07 78 04 00 08 30 
00 00 53 C0 0E 38 C3 F6 0B 93 02 70 97 0C 07 7B 
07 79 07 78 04 00 06 18 06 19 06 1A 06 1B 06 1C 
91 18 02 92 02 83 01 A0 00 00 00 00 0E 3A C0 72 
03 00 00 00 3A 56 0E 9A C0 06 0C 29 00 00 00 38 
0E 2A C0 72 01 20 00 00 00 10 38 A8 00 00 00 0C 
28 A2 2D A2 01 C0 00 00 00 00 0E AC C0 4F 02 29 
02 38 03 00 00 00 33 C0 02 A2 0C 48 00 00 00 2C 
0E 4C C0 08 02 29 0C 38 00 00 00 1C 19 40 0E 2C 
C8 71 01 30 00 00 00 10 38 28 00 00 00 0C 28 23 
27 23 01 30 00 00 00 80 26 23 01 30 00 00 00 00 
0E 23 C4 56 0C 38 00 00 00 30 01 20 00 00 00 00 
0E 32 C0 0F 02 28 82 40 0E 32 C0 05 02 29 03 00 
00 00 3B A0 01 20 00 00 00 00 0D 82 00 00 00 30 
0C 38 00 00 00 44 01 C0 00 00 00 00 0E 3C C0 08 
02 29 03 00 00 00 3B A0 0D 8C 00 00 00 44 20 20 
00 00 00 00 39 82 00 00 00 0C 03 00 00 00 3A 58 
02 2A 02 70 97 14 07 7C 07 7B 07 7A 07 79 07 78 
04 00 02 A3 02 2A 02 70 97 14 07 7C 07 7B 07 7A 
07 79 07 78 04 00 02 29 03 00 00 00 37 20 01 20 
00 00 00 10 38 A8 00 00 00 0C 28 A2 2D A2 01 C0 
00 00 00 00 0E AC C7 8C 1A 00 00 00 47 AA 02 29 
0C 38 00 00 00 10 03 00 00 00 3B A0 1A 00 00 00 
47 54 01 A0 FF FF FF FF 1A 00 00 00 47 32 91 18 
02 32 08 20 00 00 4B 34 03 00 00 00 46 C6 04 00 
06 18 06 19 06 1B 91 18 02 92 01 80 00 00 00 00 
09 80 00 00 53 C0 02 23 02 34 03 00 00 00 49 A2 
01 30 FF FF FF FF 0E 23 C0 07 02 70 97 0C 07 7B 
07 79 07 78 04 00 08 30 00 00 53 C0 0E 38 C3 F6 
0B 93 02 70 97 0C 07 7B 07 79 07 78 04 00 06 18 
06 19 06 1B 91 18 02 92 01 80 00 00 00 00 09 80 
00 00 53 C0 02 23 03 00 00 00 49 BC 01 30 FF FF 
FF FF 0E 23 C0 07 02 70 97 0C 07 7B 07 79 07 78 
04 00 08 30 00 00 53 C0 0E 38 C3 F6 0B 93 02 70 
97 0C 07 7B 07 79 07 78 04 00 06 18 06 19 06 1B 
91 18 02 92 01 80 00 00 00 00 09 80 00 00 53 C0 
02 23 02 34 02 45 03 00 00 00 49 E6 01 30 FF FF 
FF FF 0E 23 C0 07 02 70 97 0C 07 7B 07 79 07 78 
04 00 08 30 00 00 53 C0 0E 38 C3 F6 0B 93 02 70 
97 0C 07 7B 07 79 07 78 04 00 06 18 06 19 06 1B 
91 18 02 92 01 80 00 00 00 00 09 80 00 00 53 C0 
02 23 02 34 02 45 03 00 00 00 49 EE 01 30 FF FF 
FF FF 0E 23 C0 07 02 70 97 0C 07 7B 07 79 07 78 
04 00 08 30 00 00 53 C0 0E 38 C3 F6 0B 93 02 70 
97 0C 07 7B 07 79 07 78 04 00 06 18 06 19 06 1B 
91 18 08 20 00 00 53 70 01 90 FF FF FF FF 0E 29 
C0 09 01 80 00 00 53 70 19 20 98 04 0A 28 0E 29 
C7 FC 02 70 97 0C 07 7B 07 79 07 78 04 00 91 18 
04 00 01 20 00 00 20 00 0D 32 00 00 00 04 01 20 
00 00 00 00 0D 32 00 00 00 2C 04 00 01 20 00 00 
00 01 04 00 08 30 00 00 53 6C 02 43 05 42 09 40 
00 00 53 6C 02 23 04 00 30 00 00 00 00 03 04 00 
30 00 00 00 00 01 01 20 FF FF FF FF 04 00 30 00 
00 00 00 04 04 00 30 00 00 00 00 05 04 00 
@000049FE
03 00 00 00 10 DA 03 00 00 00 49 6A 04 00 
@00004A0C
03 00 00 00 10 5A 04 00 
@00004A14
48 65 6C 6C 6F 20 57 6F 72 6C 64 21 00 00 00 00 
00 00 4B 38 43 00 00 00 0A 00 00 00 
@00004B30
00 00 00 00 00 00 4B 38 00 00 00 00 00 00 4E 24 
00 00 4E 8C 00 00 4E F4 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 4A 28 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 01 33 0E AB CD 12 34 E6 6D DE EC 00 05 
00 0B 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 4F 5C 00 00 4F 5C 00 00 4F 64 
00 00 4F 64 00 00 4F 6C 00 00 4F 6C 00 00 4F 74 
00 00 4F 74 00 00 4F 7C 00 00 4F 7C 00 00 4F 84 
00 00 4F 84 00 00 4F 8C 00 00 4F 8C 00 00 4F 94 
00 00 4F 94 00 00 4F 9C 00 00 4F 9C 00 00 4F A4 
00 00 4F A4 00 00 4F AC 00 00 4F AC 00 00 4F B4 
00 00 4F B4 00 00 4F BC 00 00 4F BC 00 00 4F C4 
00 00 4F C4 00 00 4F CC 00 00 4F CC 00 00 4F D4 
00 00 4F D4 00 00 4F DC 00 00 4F DC 00 00 4F E4 
00 00 4F E4 00 00 4F EC 00 00 4F EC 00 00 4F F4 
00 00 4F F4 00 00 4F FC 00 00 4F FC 00 00 50 04 
00 00 50 04 00 00 50 0C 00 00 50 0C 00 00 50 14 
00 00 50 14 00 00 50 1C 00 00 50 1C 00 00 50 24 
00 00 50 24 00 00 50 2C 00 00 50 2C 00 00 50 34 
00 00 50 34 00 00 50 3C 00 00 50 3C 00 00 50 44 
00 00 50 44 00 00 50 4C 00 00 50 4C 00 00 50 54 
00 00 50 54 00 00 50 5C 00 00 50 5C 00 00 50 64 
00 00 50 64 00 00 50 6C 00 00 50 6C 00 00 50 74 
00 00 50 74 00 00 50 7C 00 00 50 7C 00 00 50 84 
00 00 50 84 00 00 50 8C 00 00 50 8C 00 00 50 94 
00 00 50 94 00 00 50 9C 00 00 50 9C 00 00 50 A4 
00 00 50 A4 00 00 50 AC 00 00 50 AC 00 00 50 B4 
00 00 50 B4 00 00 50 BC 00 00 50 BC 00 00 50 C4 
00 00 50 C4 00 00 50 CC 00 00 50 CC 00 00 50 D4 
00 00 50 D4 00 00 50 DC 00 00 50 DC 00 00 50 E4 
00 00 50 E4 00 00 50 EC 00 00 50 EC 00 00 50 F4 
00 00 50 F4 00 00 50 FC 00 00 50 FC 00 00 51 04 
00 00 51 04 00 00 51 0C 00 00 51 0C 00 00 51 14 
00 00 51 14 00 00 51 1C 00 00 51 1C 00 00 51 24 
00 00 51 24 00 00 51 2C 00 00 51 2C 00 00 51 34 
00 00 51 34 00 00 51 3C 00 00 51 3C 00 00 51 44 
00 00 51 44 00 00 51 4C 00 00 51 4C 00 00 51 54 
00 00 51 54 00 00 51 5C 00 00 51 5C 00 00 51 64 
00 00 51 64 00 00 51 6C 00 00 51 6C 00 00 51 74 
00 00 51 74 00 00 51 7C 00 00 51 7C 00 00 51 84 
00 00 51 84 00 00 51 8C 00 00 51 8C 00 00 51 94 
00 00 51 94 00 00 51 9C 00 00 51 9C 00 00 51 A4 
00 00 51 A4 00 00 51 AC 00 00 51 AC 00 00 51 B4 
00 00 51 B4 00 00 51 BC 00 00 51 BC 00 00 51 C4 
00 00 51 C4 00 00 51 CC 00 00 51 CC 00 00 51 D4 
00 00 51 D4 00 00 51 DC 00 00 51 DC 00 00 51 E4 
00 00 51 E4 00 00 51 EC 00 00 51 EC 00 00 51 F4 
00 00 51 F4 00 00 51 FC 00 00 51 FC 00 00 52 04 
00 00 52 04 00 00 52 0C 00 00 52 0C 00 00 52 14 
00 00 52 14 00 00 52 1C 00 00 52 1C 00 00 52 24 
00 00 52 24 00 00 52 2C 00 00 52 2C 00 00 52 34 
00 00 52 34 00 00 52 3C 00 00 52 3C 00 00 52 44 
00 00 52 44 00 00 52 4C 00 00 52 4C 00 00 52 54 
00 00 52 54 00 00 52 5C 00 00 52 5C 00 00 52 64 
00 00 52 64 00 00 52 6C 00 00 52 6C 00 00 52 74 
00 00 52 74 00 00 52 7C 00 00 52 7C 00 00 52 84 
00 00 52 84 00 00 52 8C 00 00 52 8C 00 00 52 94 
00 00 52 94 00 00 52 9C 00 00 52 9C 00 00 52 A4 
00 00 52 A4 00 00 52 AC 00 00 52 AC 00 00 52 B4 
00 00 52 B4 00 00 52 BC 00 00 52 BC 00 00 52 C4 
00 00 52 C4 00 00 52 CC 00 00 52 CC 00 00 52 D4 
00 00 52 D4 00 00 52 DC 00 00 52 DC 00 00 52 E4 
00 00 52 E4 00 00 52 EC 00 00 52 EC 00 00 52 F4 
00 00 52 F4 00 00 52 FC 00 00 52 FC 00 00 53 04 
00 00 53 04 00 00 53 0C 00 00 53 0C 00 00 53 14 
00 00 53 14 00 00 53 1C 00 00 53 1C 00 00 53 24 
00 00 53 24 00 00 53 2C 00 00 53 2C 00 00 53 34 
00 00 53 34 00 00 53 3C 00 00 53 3C 00 00 53 44 
00 00 53 44 00 00 53 4C 00 00 53 4C 00 00 53 54 
00 00 53 54 00 02 00 00 FF FF FF FF 00 00 53 C4 
@00005370
FF FF FF FF 00 00 00 00 
@00005378
FF FF FF FF 00 00 00 00 
@00005380
00 00 00 00 
